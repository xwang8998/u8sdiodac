module tap_rom(
input [1:0]oversampling_x,
input [9:0] address,
output reg signed [31:0] output_tap);

reg signed [31:0] output_1x;
reg signed [31:0] output_2x;
reg signed [31:0] output_4x;
reg signed [31:0] output_8x;

always @* begin
    if (oversampling_x==0) output_tap = output_1x[31:0];
    else if (oversampling_x==1) output_tap = output_2x[31:0];
    else if (oversampling_x==2) output_tap = output_4x[31:0];
    else output_tap = output_8x[31:0];
    end


always @* begin
    case(address)
    //10'h0: output_1x = 1073741824;
    10'h0: output_1x = 966367641;
    default: output_1x = 0;
    endcase
    end

always @* begin
    case(address)
    10'd0: output_2x = 29;
    10'd1: output_2x = 27;
    10'd2: output_2x = -89;
    10'd3: output_2x = -114;
    10'd4: output_2x = 205;
    10'd5: output_2x = 332;
    10'd6: output_2x = -395;
    10'd7: output_2x = -808;
    10'd8: output_2x = 653;
    10'd9: output_2x = 1736;
    10'd10: output_2x = -938;
    10'd11: output_2x = -3409;
    10'd12: output_2x = 1114;
    10'd13: output_2x = 6228;
    10'd14: output_2x = -915;
    10'd15: output_2x = -10722;
    10'd16: output_2x = -151;
    10'd17: output_2x = 17533;
    10'd18: output_2x = 2883;
    10'd19: output_2x = -27396;
    10'd20: output_2x = -8514;
    10'd21: output_2x = 41068;
    10'd22: output_2x = 18823;
    10'd23: output_2x = -59227;
    10'd24: output_2x = -36279;
    10'd25: output_2x = 82302;
    10'd26: output_2x = 64147;
    10'd27: output_2x = -110256;
    10'd28: output_2x = -106591;
    10'd29: output_2x = 142291;
    10'd30: output_2x = 168712;
    10'd31: output_2x = -176502;
    10'd32: output_2x = -256522;
    10'd33: output_2x = 209461;
    10'd34: output_2x = 376818;
    10'd35: output_2x = -235769;
    10'd36: output_2x = -536947;
    10'd37: output_2x = 247584;
    10'd38: output_2x = 744415;
    10'd39: output_2x = -234162;
    10'd40: output_2x = -1006369;
    10'd41: output_2x = 181437;
    10'd42: output_2x = 1328898;
    10'd43: output_2x = -71690;
    10'd44: output_2x = -1716210;
    10'd45: output_2x = -116670;
    10'd46: output_2x = 2169656;
    10'd47: output_2x = 409173;
    10'd48: output_2x = -2686663;
    10'd49: output_2x = -835183;
    10'd50: output_2x = 3259586;
    10'd51: output_2x = 1427624;
    10'd52: output_2x = -3874541;
    10'd53: output_2x = -2222547;
    10'd54: output_2x = 4510234;
    10'd55: output_2x = 3258600;
    10'd56: output_2x = -5136820;
    10'd57: output_2x = -4576492;
    10'd58: output_2x = 5714779;
    10'd59: output_2x = 6218581;
    10'd60: output_2x = -6193753;
    10'd61: output_2x = -8228841;
    10'd62: output_2x = 6511181;
    10'd63: output_2x = 10653508;
    10'd64: output_2x = -6590466;
    10'd65: output_2x = -13542926;
    10'd66: output_2x = 6338093;
    10'd67: output_2x = 16955419;
    10'd68: output_2x = -5638748;
    10'd69: output_2x = -20964582;
    10'd70: output_2x = 4346537;
    10'd71: output_2x = 25672574;
    10'd72: output_2x = -2268739;
    10'd73: output_2x = -31234575;
    10'd74: output_2x = -865491;
    10'd75: output_2x = 37905518;
    10'd76: output_2x = 5468489;
    10'd77: output_2x = -46135648;
    10'd78: output_2x = -12232426;
    10'd79: output_2x = 56786075;
    10'd80: output_2x = 22465955;
    10'd81: output_2x = -71687375;
    10'd82: output_2x = -39055800;
    10'd83: output_2x = 95413213;
    10'd84: output_2x = 69996413;
    10'd85: output_2x = -143127735;
    10'd86: output_2x = -148866205;
    10'd87: output_2x = 311192825;
    10'd88: output_2x = 846739104;
    10'd89: output_2x = 846739104;
    10'd90: output_2x = 311192825;
    10'd91: output_2x = -148866205;
    10'd92: output_2x = -143127735;
    10'd93: output_2x = 69996413;
    10'd94: output_2x = 95413213;
    10'd95: output_2x = -39055800;
    10'd96: output_2x = -71687375;
    10'd97: output_2x = 22465955;
    10'd98: output_2x = 56786075;
    10'd99: output_2x = -12232426;
    10'd100: output_2x = -46135648;
    10'd101: output_2x = 5468489;
    10'd102: output_2x = 37905518;
    10'd103: output_2x = -865491;
    10'd104: output_2x = -31234575;
    10'd105: output_2x = -2268739;
    10'd106: output_2x = 25672574;
    10'd107: output_2x = 4346537;
    10'd108: output_2x = -20964582;
    10'd109: output_2x = -5638748;
    10'd110: output_2x = 16955419;
    10'd111: output_2x = 6338093;
    10'd112: output_2x = -13542926;
    10'd113: output_2x = -6590466;
    10'd114: output_2x = 10653508;
    10'd115: output_2x = 6511181;
    10'd116: output_2x = -8228841;
    10'd117: output_2x = -6193753;
    10'd118: output_2x = 6218581;
    10'd119: output_2x = 5714779;
    10'd120: output_2x = -4576492;
    10'd121: output_2x = -5136820;
    10'd122: output_2x = 3258600;
    10'd123: output_2x = 4510234;
    10'd124: output_2x = -2222547;
    10'd125: output_2x = -3874541;
    10'd126: output_2x = 1427624;
    10'd127: output_2x = 3259586;
    10'd128: output_2x = -835183;
    10'd129: output_2x = -2686663;
    10'd130: output_2x = 409173;
    10'd131: output_2x = 2169656;
    10'd132: output_2x = -116670;
    10'd133: output_2x = -1716210;
    10'd134: output_2x = -71690;
    10'd135: output_2x = 1328898;
    10'd136: output_2x = 181437;
    10'd137: output_2x = -1006369;
    10'd138: output_2x = -234162;
    10'd139: output_2x = 744415;
    10'd140: output_2x = 247584;
    10'd141: output_2x = -536947;
    10'd142: output_2x = -235769;
    10'd143: output_2x = 376818;
    10'd144: output_2x = 209461;
    10'd145: output_2x = -256522;
    10'd146: output_2x = -176502;
    10'd147: output_2x = 168712;
    10'd148: output_2x = 142291;
    10'd149: output_2x = -106591;
    10'd150: output_2x = -110256;
    10'd151: output_2x = 64147;
    10'd152: output_2x = 82302;
    10'd153: output_2x = -36279;
    10'd154: output_2x = -59227;
    10'd155: output_2x = 18823;
    10'd156: output_2x = 41068;
    10'd157: output_2x = -8514;
    10'd158: output_2x = -27396;
    10'd159: output_2x = 2883;
    10'd160: output_2x = 17533;
    10'd161: output_2x = -151;
    10'd162: output_2x = -10722;
    10'd163: output_2x = -915;
    10'd164: output_2x = 6228;
    10'd165: output_2x = 1114;
    10'd166: output_2x = -3409;
    10'd167: output_2x = -938;
    10'd168: output_2x = 1736;
    10'd169: output_2x = 653;
    10'd170: output_2x = -808;
    10'd171: output_2x = -395;
    10'd172: output_2x = 332;
    10'd173: output_2x = 205;
    10'd174: output_2x = -114;
    10'd175: output_2x = -89;
    10'd176: output_2x = 27;
    10'd177: output_2x = 29;
    default: output_2x = 0;
    endcase
    end

always @* begin
    case(address)
    10'd0: output_4x = 22;
    10'd1: output_4x = 46;
    10'd2: output_4x = 60;
    10'd3: output_4x = 28;
    10'd4: output_4x = -67;
    10'd5: output_4x = -207;
    10'd6: output_4x = -305;
    10'd7: output_4x = -245;
    10'd8: output_4x = 53;
    10'd9: output_4x = 532;
    10'd10: output_4x = 955;
    10'd11: output_4x = 966;
    10'd12: output_4x = 296;
    10'd13: output_4x = -984;
    10'd14: output_4x = -2322;
    10'd15: output_4x = -2817;
    10'd16: output_4x = -1677;
    10'd17: output_4x = 1159;
    10'd18: output_4x = 4625;
    10'd19: output_4x = 6714;
    10'd20: output_4x = 5411;
    10'd21: output_4x = 49;
    10'd22: output_4x = -7658;
    10'd23: output_4x = -13741;
    10'd24: output_4x = -13646;
    10'd25: output_4x = -4971;
    10'd26: output_4x = 10145;
    10'd27: output_4x = 24661;
    10'd28: output_4x = 29306;
    10'd29: output_4x = 17645;
    10'd30: output_4x = -8852;
    10'd31: output_4x = -39008;
    10'd32: output_4x = -55615;
    10'd33: output_4x = -44124;
    10'd34: output_4x = -2487;
    10'd35: output_4x = 53627;
    10'd36: output_4x = 94930;
    10'd37: output_4x = 92217;
    10'd38: output_4x = 34126;
    10'd39: output_4x = -60792;
    10'd40: output_4x = -146695;
    10'd41: output_4x = -170299;
    10'd42: output_4x = -100706;
    10'd43: output_4x = 46136;
    10'd44: output_4x = 204491;
    10'd45: output_4x = 284806;
    10'd46: output_4x = 220516;
    10'd47: output_4x = 13008;
    10'd48: output_4x = -252424;
    10'd49: output_4x = -436188;
    10'd50: output_4x = -412973;
    10'd51: output_4x = -148097;
    10'd52: output_4x = 261454;
    10'd53: output_4x = 613429;
    10'd54: output_4x = 693807;
    10'd55: output_4x = 397716;
    10'd56: output_4x = -186642;
    10'd57: output_4x = -787676;
    10'd58: output_4x = -1067774;
    10'd59: output_4x = -802876;
    10'd60: output_4x = -33395;
    10'd61: output_4x = 906060;
    10'd62: output_4x = 1519225;
    10'd63: output_4x = 1398630;
    10'd64: output_4x = 473436;
    10'd65: output_4x = -887284;
    10'd66: output_4x = -2001569;
    10'd67: output_4x = -2201970;
    10'd68: output_4x = -1213820;
    10'd69: output_4x = 620817;
    10'd70: output_4x = 2427322;
    10'd71: output_4x = 3196711;
    10'd72: output_4x = 2327173;
    10'd73: output_4x = 28442;
    10'd74: output_4x = -2660989;
    10'd75: output_4x = -4317025;
    10'd76: output_4x = -3859911;
    10'd77: output_4x = -1208686;
    10'd78: output_4x = 2517186;
    10'd79: output_4x = 5431985;
    10'd80: output_4x = 5809800;
    10'd81: output_4x = 3062423;
    10'd82: output_4x = -1766067;
    10'd83: output_4x = -6333938;
    10'd84: output_4x = -8101887;
    10'd85: output_4x = -5701206;
    10'd86: output_4x = 147168;
    10'd87: output_4x = 6733251;
    10'd88: output_4x = 10565739;
    10'd89: output_4x = 9175988;
    10'd90: output_4x = 2608780;
    10'd91: output_4x = -6260902;
    10'd92: output_4x = -12916859;
    10'd93: output_4x = -13446355;
    10'd94: output_4x = -6752545;
    10'd95: output_4x = 4478160;
    10'd96: output_4x = 14743782;
    10'd97: output_4x = 18352264;
    10'd98: output_4x = 12488413;
    10'd99: output_4x = -889039;
    10'd100: output_4x = -15499160;
    10'd101: output_4x = -23591029;
    10'd102: output_4x = -19953063;
    10'd103: output_4x = -5054667;
    10'd104: output_4x = 14486653;
    10'd105: output_4x = 28699134;
    10'd106: output_4x = 29212428;
    10'd107: output_4x = 13976713;
    10'd108: output_4x = -10822018;
    10'd109: output_4x = -33030953;
    10'd110: output_4x = -40294771;
    10'd111: output_4x = -26673191;
    10'd112: output_4x = 3314848;
    10'd113: output_4x = 35708045;
    10'd114: output_4x = 53297873;
    10'd115: output_4x = 44395670;
    10'd116: output_4x = 9875005;
    10'd117: output_4x = -35459153;
    10'd118: output_4x = -68675693;
    10'd119: output_4x = -69667276;
    10'd120: output_4x = -32284737;
    10'd121: output_4x = 30071343;
    10'd122: output_4x = 88095256;
    10'd123: output_4x = 109015215;
    10'd124: output_4x = 72965206;
    10'd125: output_4x = -14138886;
    10'd126: output_4x = -117923500;
    10'd127: output_4x = -185792688;
    10'd128: output_4x = -167107657;
    10'd129: output_4x = -35492264;
    10'd130: output_4x = 196270776;
    10'd131: output_4x = 475861608;
    10'd132: output_4x = 726933705;
    10'd133: output_4x = 875216113;
    10'd134: output_4x = 875216113;
    10'd135: output_4x = 726933705;
    10'd136: output_4x = 475861608;
    10'd137: output_4x = 196270776;
    10'd138: output_4x = -35492264;
    10'd139: output_4x = -167107657;
    10'd140: output_4x = -185792688;
    10'd141: output_4x = -117923500;
    10'd142: output_4x = -14138886;
    10'd143: output_4x = 72965206;
    10'd144: output_4x = 109015215;
    10'd145: output_4x = 88095256;
    10'd146: output_4x = 30071343;
    10'd147: output_4x = -32284737;
    10'd148: output_4x = -69667276;
    10'd149: output_4x = -68675693;
    10'd150: output_4x = -35459153;
    10'd151: output_4x = 9875005;
    10'd152: output_4x = 44395670;
    10'd153: output_4x = 53297873;
    10'd154: output_4x = 35708045;
    10'd155: output_4x = 3314848;
    10'd156: output_4x = -26673191;
    10'd157: output_4x = -40294771;
    10'd158: output_4x = -33030953;
    10'd159: output_4x = -10822018;
    10'd160: output_4x = 13976713;
    10'd161: output_4x = 29212428;
    10'd162: output_4x = 28699134;
    10'd163: output_4x = 14486653;
    10'd164: output_4x = -5054667;
    10'd165: output_4x = -19953063;
    10'd166: output_4x = -23591029;
    10'd167: output_4x = -15499160;
    10'd168: output_4x = -889039;
    10'd169: output_4x = 12488413;
    10'd170: output_4x = 18352264;
    10'd171: output_4x = 14743782;
    10'd172: output_4x = 4478160;
    10'd173: output_4x = -6752545;
    10'd174: output_4x = -13446355;
    10'd175: output_4x = -12916859;
    10'd176: output_4x = -6260902;
    10'd177: output_4x = 2608780;
    10'd178: output_4x = 9175988;
    10'd179: output_4x = 10565739;
    10'd180: output_4x = 6733251;
    10'd181: output_4x = 147168;
    10'd182: output_4x = -5701206;
    10'd183: output_4x = -8101887;
    10'd184: output_4x = -6333938;
    10'd185: output_4x = -1766067;
    10'd186: output_4x = 3062423;
    10'd187: output_4x = 5809800;
    10'd188: output_4x = 5431985;
    10'd189: output_4x = 2517186;
    10'd190: output_4x = -1208686;
    10'd191: output_4x = -3859911;
    10'd192: output_4x = -4317025;
    10'd193: output_4x = -2660989;
    10'd194: output_4x = 28442;
    10'd195: output_4x = 2327173;
    10'd196: output_4x = 3196711;
    10'd197: output_4x = 2427322;
    10'd198: output_4x = 620817;
    10'd199: output_4x = -1213820;
    10'd200: output_4x = -2201970;
    10'd201: output_4x = -2001569;
    10'd202: output_4x = -887284;
    10'd203: output_4x = 473436;
    10'd204: output_4x = 1398630;
    10'd205: output_4x = 1519225;
    10'd206: output_4x = 906060;
    10'd207: output_4x = -33395;
    10'd208: output_4x = -802876;
    10'd209: output_4x = -1067774;
    10'd210: output_4x = -787676;
    10'd211: output_4x = -186642;
    10'd212: output_4x = 397716;
    10'd213: output_4x = 693807;
    10'd214: output_4x = 613429;
    10'd215: output_4x = 261454;
    10'd216: output_4x = -148097;
    10'd217: output_4x = -412973;
    10'd218: output_4x = -436188;
    10'd219: output_4x = -252424;
    10'd220: output_4x = 13008;
    10'd221: output_4x = 220516;
    10'd222: output_4x = 284806;
    10'd223: output_4x = 204491;
    10'd224: output_4x = 46136;
    10'd225: output_4x = -100706;
    10'd226: output_4x = -170299;
    10'd227: output_4x = -146695;
    10'd228: output_4x = -60792;
    10'd229: output_4x = 34126;
    10'd230: output_4x = 92217;
    10'd231: output_4x = 94930;
    10'd232: output_4x = 53627;
    10'd233: output_4x = -2487;
    10'd234: output_4x = -44124;
    10'd235: output_4x = -55615;
    10'd236: output_4x = -39008;
    10'd237: output_4x = -8852;
    10'd238: output_4x = 17645;
    10'd239: output_4x = 29306;
    10'd240: output_4x = 24661;
    10'd241: output_4x = 10145;
    10'd242: output_4x = -4971;
    10'd243: output_4x = -13646;
    10'd244: output_4x = -13741;
    10'd245: output_4x = -7658;
    10'd246: output_4x = 49;
    10'd247: output_4x = 5411;
    10'd248: output_4x = 6714;
    10'd249: output_4x = 4625;
    10'd250: output_4x = 1159;
    10'd251: output_4x = -1677;
    10'd252: output_4x = -2817;
    10'd253: output_4x = -2322;
    10'd254: output_4x = -984;
    10'd255: output_4x = 296;
    10'd256: output_4x = 966;
    10'd257: output_4x = 955;
    10'd258: output_4x = 532;
    10'd259: output_4x = 53;
    10'd260: output_4x = -245;
    10'd261: output_4x = -305;
    10'd262: output_4x = -207;
    10'd263: output_4x = -67;
    10'd264: output_4x = 28;
    10'd265: output_4x = 60;
    10'd266: output_4x = 46;
    10'd267: output_4x = 22;
    default: output_4x = 0;
    endcase
    end

always @* begin
    case(address)
    10'd0: output_8x = -19;
    10'd1: output_8x = -14;
    10'd2: output_8x = -16;
    10'd3: output_8x = -17;
    10'd4: output_8x = -13;
    10'd5: output_8x = -7;
    10'd6: output_8x = 2;
    10'd7: output_8x = 16;
    10'd8: output_8x = 30;
    10'd9: output_8x = 45;
    10'd10: output_8x = 55;
    10'd11: output_8x = 62;
    10'd12: output_8x = 59;
    10'd13: output_8x = 47;
    10'd14: output_8x = 27;
    10'd15: output_8x = -1;
    10'd16: output_8x = -36;
    10'd17: output_8x = -72;
    10'd18: output_8x = -104;
    10'd19: output_8x = -125;
    10'd20: output_8x = -131;
    10'd21: output_8x = -117;
    10'd22: output_8x = -83;
    10'd23: output_8x = -30;
    10'd24: output_8x = 36;
    10'd25: output_8x = 110;
    10'd26: output_8x = 181;
    10'd27: output_8x = 236;
    10'd28: output_8x = 265;
    10'd29: output_8x = 259;
    10'd30: output_8x = 213;
    10'd31: output_8x = 127;
    10'd32: output_8x = 9;
    10'd33: output_8x = -126;
    10'd34: output_8x = -267;
    10'd35: output_8x = -387;
    10'd36: output_8x = -469;
    10'd37: output_8x = -493;
    10'd38: output_8x = -446;
    10'd39: output_8x = -326;
    10'd40: output_8x = -141;
    10'd41: output_8x = 90;
    10'd42: output_8x = 342;
    10'd43: output_8x = 576;
    10'd44: output_8x = 758;
    10'd45: output_8x = 853;
    10'd46: output_8x = 834;
    10'd47: output_8x = 690;
    10'd48: output_8x = 424;
    10'd49: output_8x = 63;
    10'd50: output_8x = -352;
    10'd51: output_8x = -770;
    10'd52: output_8x = -1126;
    10'd53: output_8x = -1362;
    10'd54: output_8x = -1427;
    10'd55: output_8x = -1290;
    10'd56: output_8x = -948;
    10'd57: output_8x = -427;
    10'd58: output_8x = 216;
    10'd59: output_8x = 906;
    10'd60: output_8x = 1543;
    10'd61: output_8x = 2028;
    10'd62: output_8x = 2273;
    10'd63: output_8x = 2214;
    10'd64: output_8x = 1826;
    10'd65: output_8x = 1128;
    10'd66: output_8x = 190;
    10'd67: output_8x = -877;
    10'd68: output_8x = -1934;
    10'd69: output_8x = -2824;
    10'd70: output_8x = -3399;
    10'd71: output_8x = -3542;
    10'd72: output_8x = -3186;
    10'd73: output_8x = -2331;
    10'd74: output_8x = -1049;
    10'd75: output_8x = 514;
    10'd76: output_8x = 2165;
    10'd77: output_8x = 3670;
    10'd78: output_8x = 4794;
    10'd79: output_8x = 5338;
    10'd80: output_8x = 5165;
    10'd81: output_8x = 4228;
    10'd82: output_8x = 2589;
    10'd83: output_8x = 417;
    10'd84: output_8x = -2023;
    10'd85: output_8x = -4406;
    10'd86: output_8x = -6381;
    10'd87: output_8x = -7623;
    10'd88: output_8x = -7884;
    10'd89: output_8x = -7033;
    10'd90: output_8x = -5091;
    10'd91: output_8x = -2238;
    10'd92: output_8x = 1197;
    10'd93: output_8x = 4773;
    10'd94: output_8x = 7987;
    10'd95: output_8x = 10341;
    10'd96: output_8x = 11419;
    10'd97: output_8x = 10953;
    10'd98: output_8x = 8873;
    10'd99: output_8x = 5337;
    10'd100: output_8x = 729;
    10'd101: output_8x = -4382;
    10'd102: output_8x = -9305;
    10'd103: output_8x = -13314;
    10'd104: output_8x = -15757;
    10'd105: output_8x = -16148;
    10'd106: output_8x = -14260;
    10'd107: output_8x = -10172;
    10'd108: output_8x = -4289;
    10'd109: output_8x = 2692;
    10'd110: output_8x = 9862;
    10'd111: output_8x = 16206;
    10'd112: output_8x = 20748;
    10'd113: output_8x = 22690;
    10'd114: output_8x = 21546;
    10'd115: output_8x = 17232;
    10'd116: output_8x = 10114;
    10'd117: output_8x = 990;
    10'd118: output_8x = -8989;
    10'd119: output_8x = -18466;
    10'd120: output_8x = -26043;
    10'd121: output_8x = -30490;
    10'd122: output_8x = -30930;
    10'd123: output_8x = -26993;
    10'd124: output_8x = -18909;
    10'd125: output_8x = -7520;
    10'd126: output_8x = 5796;
    10'd127: output_8x = 19284;
    10'd128: output_8x = 31029;
    10'd129: output_8x = 39225;
    10'd130: output_8x = 42440;
    10'd131: output_8x = 39850;
    10'd132: output_8x = 31401;
    10'd133: output_8x = 17871;
    10'd134: output_8x = 823;
    10'd135: output_8x = -17565;
    10'd136: output_8x = -34770;
    10'd137: output_8x = -48256;
    10'd138: output_8x = -55837;
    10'd139: output_8x = -56017;
    10'd140: output_8x = -48252;
    10'd141: output_8x = -33092;
    10'd142: output_8x = -12180;
    10'd143: output_8x = 11902;
    10'd144: output_8x = 35951;
    10'd145: output_8x = 56541;
    10'd146: output_8x = 70508;
    10'd147: output_8x = 75418;
    10'd148: output_8x = 69959;
    10'd149: output_8x = 54213;
    10'd150: output_8x = 29727;
    10'd151: output_8x = -596;
    10'd152: output_8x = -32843;
    10'd153: output_8x = -62558;
    10'd154: output_8x = -85354;
    10'd155: output_8x = -97544;
    10'd156: output_8x = -96708;
    10'd157: output_8x = -82121;
    10'd158: output_8x = -54967;
    10'd159: output_8x = -18292;
    10'd160: output_8x = 23307;
    10'd161: output_8x = 64249;
    10'd162: output_8x = 98684;
    10'd163: output_8x = 121320;
    10'd164: output_8x = 128211;
    10'd165: output_8x = 117396;
    10'd166: output_8x = 89308;
    10'd167: output_8x = 46858;
    10'd168: output_8x = -4825;
    10'd169: output_8x = -58992;
    10'd170: output_8x = -108121;
    10'd171: output_8x = -144952;
    10'd172: output_8x = -163527;
    10'd173: output_8x = -160118;
    10'd174: output_8x = -133887;
    10'd175: output_8x = -87184;
    10'd176: output_8x = -25398;
    10'd177: output_8x = 43625;
    10'd178: output_8x = 110553;
    10'd179: output_8x = 165798;
    10'd180: output_8x = 200869;
    10'd181: output_8x = 209632;
    10'd182: output_8x = 189325;
    10'd183: output_8x = 141140;
    10'd184: output_8x = 70283;
    10'd185: output_8x = -14531;
    10'd186: output_8x = -102123;
    10'd187: output_8x = -180279;
    10'd188: output_8x = -237428;
    10'd189: output_8x = -264320;
    10'd190: output_8x = -255464;
    10'd191: output_8x = -210114;
    10'd192: output_8x = -132643;
    10'd193: output_8x = -32205;
    10'd194: output_8x = 78294;
    10'd195: output_8x = 183823;
    10'd196: output_8x = 269223;
    10'd197: output_8x = 321354;
    10'd198: output_8x = 331064;
    10'd199: output_8x = 294688;
    10'd200: output_8x = 214880;
    10'd201: output_8x = 100561;
    10'd202: output_8x = -33996;
    10'd203: output_8x = -170910;
    10'd204: output_8x = -291011;
    10'd205: output_8x = -376494;
    10'd206: output_8x = -413499;
    10'd207: output_8x = -394281;
    10'd208: output_8x = -318616;
    10'd209: output_8x = -194231;
    10'd210: output_8x = -36122;
    10'd211: output_8x = 135189;
    10'd212: output_8x = 296265;
    10'd213: output_8x = 423915;
    10'd214: output_8x = 498473;
    10'd215: output_8x = 506758;
    10'd216: output_8x = 444261;
    10'd217: output_8x = 316214;
    10'd218: output_8x = 137346;
    10'd219: output_8x = -69720;
    10'd220: output_8x = -277269;
    10'd221: output_8x = -456139;
    10'd222: output_8x = -579769;
    10'd223: output_8x = -628064;
    10'd224: output_8x = -590549;
    10'd225: output_8x = -468315;
    10'd226: output_8x = -274425;
    10'd227: output_8x = -32656;
    10'd228: output_8x = 225326;
    10'd229: output_8x = 464062;
    10'd230: output_8x = 649093;
    10'd231: output_8x = 751870;
    10'd232: output_8x = 754056;
    10'd233: output_8x = 650584;
    10'd234: output_8x = 451005;
    10'd235: output_8x = 178829;
    10'd236: output_8x = -131131;
    10'd237: output_8x = -437129;
    10'd238: output_8x = -696031;
    10'd239: output_8x = -869323;
    10'd240: output_8x = -928744;
    10'd241: output_8x = -860726;
    10'd242: output_8x = -668984;
    10'd243: output_8x = -374776;
    10'd244: output_8x = -14717;
    10'd245: output_8x = 363669;
    10'd246: output_8x = 708147;
    10'd247: output_8x = 968884;
    10'd248: output_8x = 1105573;
    10'd249: output_8x = 1093517;
    10'd250: output_8x = 927795;
    10'd251: output_8x = 624835;
    10'd252: output_8x = 221044;
    10'd253: output_8x = -231417;
    10'd254: output_8x = -671277;
    10'd255: output_8x = -1036349;
    10'd256: output_8x = -1272228;
    10'd257: output_8x = -1340267;
    10'd258: output_8x = -1223685;
    10'd259: output_8x = -930866;
    10'd260: output_8x = -495263;
    10'd261: output_8x = 28220;
    10'd262: output_8x = 570022;
    10'd263: output_8x = 1055052;
    10'd264: output_8x = 1413000;
    10'd265: output_8x = 1588394;
    10'd266: output_8x = 1549012;
    10'd267: output_8x = 1291374;
    10'd268: output_8x = 842436;
    10'd269: output_8x = 257069;
    10'd270: output_8x = -388457;
    10'd271: output_8x = -1006304;
    10'd272: output_8x = -1508881;
    10'd273: output_8x = -1821147;
    10'd274: output_8x = -1891635;
    10'd275: output_8x = -1700631;
    10'd276: output_8x = -1264235;
    10'd277: output_8x = -633546;
    10'd278: output_8x = 111070;
    10'd279: output_8x = 870071;
    10'd280: output_8x = 1537900;
    10'd281: output_8x = 2017541;
    10'd282: output_8x = 2234444;
    10'd283: output_8x = 2147859;
    10'd284: output_8x = 1757880;
    10'd285: output_8x = 1107056;
    10'd286: output_8x = 276095;
    10'd287: output_8x = -625930;
    10'd288: output_8x = -1475743;
    10'd289: output_8x = -2152565;
    10'd290: output_8x = -2555112;
    10'd291: output_8x = -2616534;
    10'd292: output_8x = -2315094;
    10'd293: output_8x = -1678950;
    10'd294: output_8x = -784133;
    10'd295: output_8x = 254257;
    10'd296: output_8x = 1296666;
    10'd297: output_8x = 2197669;
    10'd298: output_8x = 2826096;
    10'd299: output_8x = 3083906;
    10'd300: output_8x = 2921160;
    10'd301: output_8x = 2344802;
    10'd302: output_8x = 1419823;
    10'd303: output_8x = 262349;
    10'd304: output_8x = -974698;
    10'd305: output_8x = -2121604;
    10'd306: output_8x = -3014965;
    10'd307: output_8x = -3520761;
    10'd308: output_8x = -3554164;
    10'd309: output_8x = -3093203;
    10'd310: output_8x = -2184137;
    10'd311: output_8x = -937472;
    10'd312: output_8x = 485126;
    10'd313: output_8x = 1891572;
    10'd314: output_8x = 3085086;
    10'd315: output_8x = 3891515;
    10'd316: output_8x = 4184469;
    10'd317: output_8x = 3904694;
    10'd318: output_8x = 3070739;
    10'd319: output_8x = 1779156;
    10'd320: output_8x = 193788;
    10'd321: output_8x = -1474717;
    10'd322: output_8x = -2996660;
    10'd323: output_8x = -4154679;
    10'd324: output_8x = -4774526;
    10'd325: output_8x = -4750912;
    10'd326: output_8x = -4064614;
    10'd327: output_8x = -2788162;
    10'd328: output_8x = -1078927;
    10'd329: output_8x = 839895;
    10'd330: output_8x = 2708145;
    10'd331: output_8x = 4263710;
    10'd332: output_8x = 5279038;
    10'd333: output_8x = 5594061;
    10'd334: output_8x = 5140851;
    10'd335: output_8x = 3956251;
    10'd336: output_8x = 2180322;
    10'd337: output_8x = 40327;
    10'd338: output_8x = -2177990;
    10'd339: output_8x = -4168267;
    10'd340: output_8x = -5645541;
    10'd341: output_8x = -6386711;
    10'd342: output_8x = -6263725;
    10'd343: output_8x = -5264637;
    10'd344: output_8x = -3499173;
    10'd345: output_8x = -1187522;
    10'd346: output_8x = 1366667;
    10'd347: output_8x = 3815816;
    10'd348: output_8x = 5815392;
    10'd349: output_8x = 7072026;
    10'd350: output_8x = 7386093;
    10'd351: output_8x = 6682642;
    10'd352: output_8x = 5025954;
    10'd353: output_8x = 2615196;
    10'd354: output_8x = -238880;
    10'd355: output_8x = -3153567;
    10'd356: output_8x = -5725133;
    10'd357: output_8x = -7584377;
    10'd358: output_8x = -8449188;
    10'd359: output_8x = -8166678;
    10'd360: output_8x = -6738701;
    10'd361: output_8x = -4326639;
    10'd362: output_8x = -1234125;
    10'd363: output_8x = 2130608;
    10'd364: output_8x = 5308178;
    10'd365: output_8x = 7850343;
    10'd366: output_8x = 9382776;
    10'd367: output_8x = 9659561;
    10'd368: output_8x = 8601586;
    10'd369: output_8x = 6312932;
    10'd370: output_8x = 3072302;
    10'd371: output_8x = -700143;
    10'd372: output_8x = -4496708;
    10'd373: output_8x = -7789999;
    10'd374: output_8x = -10105681;
    10'd375: output_8x = -11090189;
    10'd376: output_8x = -10563801;
    10'd377: output_8x = -8551218;
    10'd378: output_8x = -5284687;
    10'd379: output_8x = -1178336;
    10'd380: output_8x = 3223604;
    10'd381: output_8x = 7318351;
    10'd382: output_8x = 10526528;
    10'd383: output_8x = 12373509;
    10'd384: output_8x = 12558782;
    10'd385: output_8x = 11003312;
    10'd386: output_8x = 7867624;
    10'd387: output_8x = 3537140;
    10'd388: output_8x = -1424211;
    10'd389: output_8x = -6346701;
    10'd390: output_8x = -10544528;
    10'd391: output_8x = -13410647;
    10'd392: output_8x = -14503698;
    10'd393: output_8x = -13614667;
    10'd394: output_8x = -10803404;
    10'd395: output_8x = -6398933;
    10'd396: output_8x = -962368;
    10'd397: output_8x = 4783606;
    10'd398: output_8x = 10049979;
    10'd399: output_8x = 14088922;
    10'd400: output_8x = 16299041;
    10'd401: output_8x = 16313686;
    10'd402: output_8x = 14059485;
    10'd403: output_8x = 9776052;
    10'd404: output_8x = 3992850;
    10'd405: output_8x = -2534940;
    10'd406: output_8x = -8923980;
    10'd407: output_8x = -14281293;
    10'd408: output_8x = -17827996;
    10'd409: output_8x = -19011228;
    10'd410: output_8x = -17588359;
    10'd411: output_8x = -13670915;
    10'd412: output_8x = -7720777;
    10'd413: output_8x = -497652;
    10'd414: output_8x = 7036537;
    10'd415: output_8x = 13844478;
    10'd416: output_8x = 18954973;
    10'd417: output_8x = 21599993;
    10'd418: output_8x = 21328140;
    10'd419: output_8x = 18077993;
    10'd420: output_8x = 12199852;
    10'd421: output_8x = 4421129;
    10'd422: output_8x = -4241738;
    10'd423: output_8x = -12614431;
    10'd424: output_8x = -19522269;
    10'd425: output_8x = -23953202;
    10'd426: output_8x = -25203895;
    10'd427: output_8x = -22988094;
    10'd428: output_8x = -17490995;
    10'd429: output_8x = -9360207;
    10'd430: output_8x = 367655;
    10'd431: output_8x = 10396858;
    10'd432: output_8x = 19342923;
    10'd433: output_8x = 25921422;
    10'd434: output_8x = 29129705;
    10'd435: output_8x = 28396244;
    10'd436: output_8x = 23675761;
    10'd437: output_8x = 15475051;
    10'd438: output_8x = 4803394;
    10'd439: output_8x = -6948371;
    10'd440: output_8x = -18186085;
    10'd441: output_8x = -27325347;
    10'd442: output_8x = -33011387;
    10'd443: output_8x = -34315670;
    10'd444: output_8x = -30881251;
    10'd445: output_8x = -22994877;
    10'd446: output_8x = -11573068;
    10'd447: output_8x = 1939275;
    10'd448: output_8x = 15747264;
    10'd449: output_8x = 27939933;
    10'd450: output_8x = 36749772;
    10'd451: output_8x = 40803261;
    10'd452: output_8x = 39327625;
    10'd453: output_8x = 32283642;
    10'd454: output_8x = 20403141;
    10'd455: output_8x = 5122049;
    10'd456: output_8x = -11586353;
    10'd457: output_8x = -27459480;
    10'd458: output_8x = -40244410;
    10'd459: output_8x = -48009229;
    10'd460: output_8x = -49424743;
    10'd461: output_8x = -43976818;
    10'd462: output_8x = -32077170;
    10'd463: output_8x = -15052768;
    10'd464: output_8x = 4990471;
    10'd465: output_8x = 25417265;
    10'd466: output_8x = 43397500;
    10'd467: output_8x = 56284639;
    10'd468: output_8x = 61989041;
    10'd469: output_8x = 59295528;
    10'd470: output_8x = 48079494;
    10'd471: output_8x = 29387144;
    10'd472: output_8x = 5361761;
    10'd473: output_8x = -20982545;
    10'd474: output_8x = -46117878;
    10'd475: output_8x = -66450236;
    10'd476: output_8x = -78803650;
    10'd477: output_8x = -80878864;
    10'd478: output_8x = -71624595;
    10'd479: output_8x = -51467368;
    10'd480: output_8x = -22361203;
    10'd481: output_8x = 12360575;
    10'd482: output_8x = 48324848;
    10'd483: output_8x = 80618256;
    10'd484: output_8x = 104393673;
    10'd485: output_8x = 115514007;
    10'd486: output_8x = 111155346;
    10'd487: output_8x = 90292157;
    10'd488: output_8x = 53997556;
    10'd489: output_8x = 5510631;
    10'd490: output_8x = -49951638;
    10'd491: output_8x = -105630862;
    10'd492: output_8x = -153875285;
    10'd493: output_8x = -186935969;
    10'd494: output_8x = -197827466;
    10'd495: output_8x = -181158231;
    10'd496: output_8x = -133835661;
    10'd497: output_8x = -55561196;
    10'd498: output_8x = 50948326;
    10'd499: output_8x = 180048300;
    10'd500: output_8x = 323564692;
    10'd501: output_8x = 471470497;
    10'd502: output_8x = 612776116;
    10'd503: output_8x = 736544613;
    10'd504: output_8x = 832927451;
    10'd505: output_8x = 894112424;
    10'd506: output_8x = 915083602;
    10'd507: output_8x = 894112424;
    10'd508: output_8x = 832927451;
    10'd509: output_8x = 736544613;
    10'd510: output_8x = 612776116;
    10'd511: output_8x = 471470497;
    10'd512: output_8x = 323564692;
    10'd513: output_8x = 180048300;
    10'd514: output_8x = 50948326;
    10'd515: output_8x = -55561196;
    10'd516: output_8x = -133835661;
    10'd517: output_8x = -181158231;
    10'd518: output_8x = -197827466;
    10'd519: output_8x = -186935969;
    10'd520: output_8x = -153875285;
    10'd521: output_8x = -105630862;
    10'd522: output_8x = -49951638;
    10'd523: output_8x = 5510631;
    10'd524: output_8x = 53997556;
    10'd525: output_8x = 90292157;
    10'd526: output_8x = 111155346;
    10'd527: output_8x = 115514007;
    10'd528: output_8x = 104393673;
    10'd529: output_8x = 80618256;
    10'd530: output_8x = 48324848;
    10'd531: output_8x = 12360575;
    10'd532: output_8x = -22361203;
    10'd533: output_8x = -51467368;
    10'd534: output_8x = -71624595;
    10'd535: output_8x = -80878864;
    10'd536: output_8x = -78803650;
    10'd537: output_8x = -66450236;
    10'd538: output_8x = -46117878;
    10'd539: output_8x = -20982545;
    10'd540: output_8x = 5361761;
    10'd541: output_8x = 29387144;
    10'd542: output_8x = 48079494;
    10'd543: output_8x = 59295528;
    10'd544: output_8x = 61989041;
    10'd545: output_8x = 56284639;
    10'd546: output_8x = 43397500;
    10'd547: output_8x = 25417265;
    10'd548: output_8x = 4990471;
    10'd549: output_8x = -15052768;
    10'd550: output_8x = -32077170;
    10'd551: output_8x = -43976818;
    10'd552: output_8x = -49424743;
    10'd553: output_8x = -48009229;
    10'd554: output_8x = -40244410;
    10'd555: output_8x = -27459480;
    10'd556: output_8x = -11586353;
    10'd557: output_8x = 5122049;
    10'd558: output_8x = 20403141;
    10'd559: output_8x = 32283642;
    10'd560: output_8x = 39327625;
    10'd561: output_8x = 40803261;
    10'd562: output_8x = 36749772;
    10'd563: output_8x = 27939933;
    10'd564: output_8x = 15747264;
    10'd565: output_8x = 1939275;
    10'd566: output_8x = -11573068;
    10'd567: output_8x = -22994877;
    10'd568: output_8x = -30881251;
    10'd569: output_8x = -34315670;
    10'd570: output_8x = -33011387;
    10'd571: output_8x = -27325347;
    10'd572: output_8x = -18186085;
    10'd573: output_8x = -6948371;
    10'd574: output_8x = 4803394;
    10'd575: output_8x = 15475051;
    10'd576: output_8x = 23675761;
    10'd577: output_8x = 28396244;
    10'd578: output_8x = 29129705;
    10'd579: output_8x = 25921422;
    10'd580: output_8x = 19342923;
    10'd581: output_8x = 10396858;
    10'd582: output_8x = 367655;
    10'd583: output_8x = -9360207;
    10'd584: output_8x = -17490995;
    10'd585: output_8x = -22988094;
    10'd586: output_8x = -25203895;
    10'd587: output_8x = -23953202;
    10'd588: output_8x = -19522269;
    10'd589: output_8x = -12614431;
    10'd590: output_8x = -4241738;
    10'd591: output_8x = 4421129;
    10'd592: output_8x = 12199852;
    10'd593: output_8x = 18077993;
    10'd594: output_8x = 21328140;
    10'd595: output_8x = 21599993;
    10'd596: output_8x = 18954973;
    10'd597: output_8x = 13844478;
    10'd598: output_8x = 7036537;
    10'd599: output_8x = -497652;
    10'd600: output_8x = -7720777;
    10'd601: output_8x = -13670915;
    10'd602: output_8x = -17588359;
    10'd603: output_8x = -19011228;
    10'd604: output_8x = -17827996;
    10'd605: output_8x = -14281293;
    10'd606: output_8x = -8923980;
    10'd607: output_8x = -2534940;
    10'd608: output_8x = 3992850;
    10'd609: output_8x = 9776052;
    10'd610: output_8x = 14059485;
    10'd611: output_8x = 16313686;
    10'd612: output_8x = 16299041;
    10'd613: output_8x = 14088922;
    10'd614: output_8x = 10049979;
    10'd615: output_8x = 4783606;
    10'd616: output_8x = -962368;
    10'd617: output_8x = -6398933;
    10'd618: output_8x = -10803404;
    10'd619: output_8x = -13614667;
    10'd620: output_8x = -14503698;
    10'd621: output_8x = -13410647;
    10'd622: output_8x = -10544528;
    10'd623: output_8x = -6346701;
    10'd624: output_8x = -1424211;
    10'd625: output_8x = 3537140;
    10'd626: output_8x = 7867624;
    10'd627: output_8x = 11003312;
    10'd628: output_8x = 12558782;
    10'd629: output_8x = 12373509;
    10'd630: output_8x = 10526528;
    10'd631: output_8x = 7318351;
    10'd632: output_8x = 3223604;
    10'd633: output_8x = -1178336;
    10'd634: output_8x = -5284687;
    10'd635: output_8x = -8551218;
    10'd636: output_8x = -10563801;
    10'd637: output_8x = -11090189;
    10'd638: output_8x = -10105681;
    10'd639: output_8x = -7789999;
    10'd640: output_8x = -4496708;
    10'd641: output_8x = -700143;
    10'd642: output_8x = 3072302;
    10'd643: output_8x = 6312932;
    10'd644: output_8x = 8601586;
    10'd645: output_8x = 9659561;
    10'd646: output_8x = 9382776;
    10'd647: output_8x = 7850343;
    10'd648: output_8x = 5308178;
    10'd649: output_8x = 2130608;
    10'd650: output_8x = -1234125;
    10'd651: output_8x = -4326639;
    10'd652: output_8x = -6738701;
    10'd653: output_8x = -8166678;
    10'd654: output_8x = -8449188;
    10'd655: output_8x = -7584377;
    10'd656: output_8x = -5725133;
    10'd657: output_8x = -3153567;
    10'd658: output_8x = -238880;
    10'd659: output_8x = 2615196;
    10'd660: output_8x = 5025954;
    10'd661: output_8x = 6682642;
    10'd662: output_8x = 7386093;
    10'd663: output_8x = 7072026;
    10'd664: output_8x = 5815392;
    10'd665: output_8x = 3815816;
    10'd666: output_8x = 1366667;
    10'd667: output_8x = -1187522;
    10'd668: output_8x = -3499173;
    10'd669: output_8x = -5264637;
    10'd670: output_8x = -6263725;
    10'd671: output_8x = -6386711;
    10'd672: output_8x = -5645541;
    10'd673: output_8x = -4168267;
    10'd674: output_8x = -2177990;
    10'd675: output_8x = 40327;
    10'd676: output_8x = 2180322;
    10'd677: output_8x = 3956251;
    10'd678: output_8x = 5140851;
    10'd679: output_8x = 5594061;
    10'd680: output_8x = 5279038;
    10'd681: output_8x = 4263710;
    10'd682: output_8x = 2708145;
    10'd683: output_8x = 839895;
    10'd684: output_8x = -1078927;
    10'd685: output_8x = -2788162;
    10'd686: output_8x = -4064614;
    10'd687: output_8x = -4750912;
    10'd688: output_8x = -4774526;
    10'd689: output_8x = -4154679;
    10'd690: output_8x = -2996660;
    10'd691: output_8x = -1474717;
    10'd692: output_8x = 193788;
    10'd693: output_8x = 1779156;
    10'd694: output_8x = 3070739;
    10'd695: output_8x = 3904694;
    10'd696: output_8x = 4184469;
    10'd697: output_8x = 3891515;
    10'd698: output_8x = 3085086;
    10'd699: output_8x = 1891572;
    10'd700: output_8x = 485126;
    10'd701: output_8x = -937472;
    10'd702: output_8x = -2184137;
    10'd703: output_8x = -3093203;
    10'd704: output_8x = -3554164;
    10'd705: output_8x = -3520761;
    10'd706: output_8x = -3014965;
    10'd707: output_8x = -2121604;
    10'd708: output_8x = -974698;
    10'd709: output_8x = 262349;
    10'd710: output_8x = 1419823;
    10'd711: output_8x = 2344802;
    10'd712: output_8x = 2921160;
    10'd713: output_8x = 3083906;
    10'd714: output_8x = 2826096;
    10'd715: output_8x = 2197669;
    10'd716: output_8x = 1296666;
    10'd717: output_8x = 254257;
    10'd718: output_8x = -784133;
    10'd719: output_8x = -1678950;
    10'd720: output_8x = -2315094;
    10'd721: output_8x = -2616534;
    10'd722: output_8x = -2555112;
    10'd723: output_8x = -2152565;
    10'd724: output_8x = -1475743;
    10'd725: output_8x = -625930;
    10'd726: output_8x = 276095;
    10'd727: output_8x = 1107056;
    10'd728: output_8x = 1757880;
    10'd729: output_8x = 2147859;
    10'd730: output_8x = 2234444;
    10'd731: output_8x = 2017541;
    10'd732: output_8x = 1537900;
    10'd733: output_8x = 870071;
    10'd734: output_8x = 111070;
    10'd735: output_8x = -633546;
    10'd736: output_8x = -1264235;
    10'd737: output_8x = -1700631;
    10'd738: output_8x = -1891635;
    10'd739: output_8x = -1821147;
    10'd740: output_8x = -1508881;
    10'd741: output_8x = -1006304;
    10'd742: output_8x = -388457;
    10'd743: output_8x = 257069;
    10'd744: output_8x = 842436;
    10'd745: output_8x = 1291374;
    10'd746: output_8x = 1549012;
    10'd747: output_8x = 1588394;
    10'd748: output_8x = 1413000;
    10'd749: output_8x = 1055052;
    10'd750: output_8x = 570022;
    10'd751: output_8x = 28220;
    10'd752: output_8x = -495263;
    10'd753: output_8x = -930866;
    10'd754: output_8x = -1223685;
    10'd755: output_8x = -1340267;
    10'd756: output_8x = -1272228;
    10'd757: output_8x = -1036349;
    10'd758: output_8x = -671277;
    10'd759: output_8x = -231417;
    10'd760: output_8x = 221044;
    10'd761: output_8x = 624835;
    10'd762: output_8x = 927795;
    10'd763: output_8x = 1093517;
    10'd764: output_8x = 1105573;
    10'd765: output_8x = 968884;
    10'd766: output_8x = 708147;
    10'd767: output_8x = 363669;
    10'd768: output_8x = -14717;
    10'd769: output_8x = -374776;
    10'd770: output_8x = -668984;
    10'd771: output_8x = -860726;
    10'd772: output_8x = -928744;
    10'd773: output_8x = -869323;
    10'd774: output_8x = -696031;
    10'd775: output_8x = -437129;
    10'd776: output_8x = -131131;
    10'd777: output_8x = 178829;
    10'd778: output_8x = 451005;
    10'd779: output_8x = 650584;
    10'd780: output_8x = 754056;
    10'd781: output_8x = 751870;
    10'd782: output_8x = 649093;
    10'd783: output_8x = 464062;
    10'd784: output_8x = 225326;
    10'd785: output_8x = -32656;
    10'd786: output_8x = -274425;
    10'd787: output_8x = -468315;
    10'd788: output_8x = -590549;
    10'd789: output_8x = -628064;
    10'd790: output_8x = -579769;
    10'd791: output_8x = -456139;
    10'd792: output_8x = -277269;
    10'd793: output_8x = -69720;
    10'd794: output_8x = 137346;
    10'd795: output_8x = 316214;
    10'd796: output_8x = 444261;
    10'd797: output_8x = 506758;
    10'd798: output_8x = 498473;
    10'd799: output_8x = 423915;
    10'd800: output_8x = 296265;
    10'd801: output_8x = 135189;
    10'd802: output_8x = -36122;
    10'd803: output_8x = -194231;
    10'd804: output_8x = -318616;
    10'd805: output_8x = -394281;
    10'd806: output_8x = -413499;
    10'd807: output_8x = -376494;
    10'd808: output_8x = -291011;
    10'd809: output_8x = -170910;
    10'd810: output_8x = -33996;
    10'd811: output_8x = 100561;
    10'd812: output_8x = 214880;
    10'd813: output_8x = 294688;
    10'd814: output_8x = 331064;
    10'd815: output_8x = 321354;
    10'd816: output_8x = 269223;
    10'd817: output_8x = 183823;
    10'd818: output_8x = 78294;
    10'd819: output_8x = -32205;
    10'd820: output_8x = -132643;
    10'd821: output_8x = -210114;
    10'd822: output_8x = -255464;
    10'd823: output_8x = -264320;
    10'd824: output_8x = -237428;
    10'd825: output_8x = -180279;
    10'd826: output_8x = -102123;
    10'd827: output_8x = -14531;
    10'd828: output_8x = 70283;
    10'd829: output_8x = 141140;
    10'd830: output_8x = 189325;
    10'd831: output_8x = 209632;
    10'd832: output_8x = 200869;
    10'd833: output_8x = 165798;
    10'd834: output_8x = 110553;
    10'd835: output_8x = 43625;
    10'd836: output_8x = -25398;
    10'd837: output_8x = -87184;
    10'd838: output_8x = -133887;
    10'd839: output_8x = -160118;
    10'd840: output_8x = -163527;
    10'd841: output_8x = -144952;
    10'd842: output_8x = -108121;
    10'd843: output_8x = -58992;
    10'd844: output_8x = -4825;
    10'd845: output_8x = 46858;
    10'd846: output_8x = 89308;
    10'd847: output_8x = 117396;
    10'd848: output_8x = 128211;
    10'd849: output_8x = 121320;
    10'd850: output_8x = 98684;
    10'd851: output_8x = 64249;
    10'd852: output_8x = 23307;
    10'd853: output_8x = -18292;
    10'd854: output_8x = -54967;
    10'd855: output_8x = -82121;
    10'd856: output_8x = -96708;
    10'd857: output_8x = -97544;
    10'd858: output_8x = -85354;
    10'd859: output_8x = -62558;
    10'd860: output_8x = -32843;
    10'd861: output_8x = -596;
    10'd862: output_8x = 29727;
    10'd863: output_8x = 54213;
    10'd864: output_8x = 69959;
    10'd865: output_8x = 75418;
    10'd866: output_8x = 70508;
    10'd867: output_8x = 56541;
    10'd868: output_8x = 35951;
    10'd869: output_8x = 11902;
    10'd870: output_8x = -12180;
    10'd871: output_8x = -33092;
    10'd872: output_8x = -48252;
    10'd873: output_8x = -56017;
    10'd874: output_8x = -55837;
    10'd875: output_8x = -48256;
    10'd876: output_8x = -34770;
    10'd877: output_8x = -17565;
    10'd878: output_8x = 823;
    10'd879: output_8x = 17871;
    10'd880: output_8x = 31401;
    10'd881: output_8x = 39850;
    10'd882: output_8x = 42440;
    10'd883: output_8x = 39225;
    10'd884: output_8x = 31029;
    10'd885: output_8x = 19284;
    10'd886: output_8x = 5796;
    10'd887: output_8x = -7520;
    10'd888: output_8x = -18909;
    10'd889: output_8x = -26993;
    10'd890: output_8x = -30930;
    10'd891: output_8x = -30490;
    10'd892: output_8x = -26043;
    10'd893: output_8x = -18466;
    10'd894: output_8x = -8989;
    10'd895: output_8x = 990;
    10'd896: output_8x = 10114;
    10'd897: output_8x = 17232;
    10'd898: output_8x = 21546;
    10'd899: output_8x = 22690;
    10'd900: output_8x = 20748;
    10'd901: output_8x = 16206;
    10'd902: output_8x = 9862;
    10'd903: output_8x = 2692;
    10'd904: output_8x = -4289;
    10'd905: output_8x = -10172;
    10'd906: output_8x = -14260;
    10'd907: output_8x = -16148;
    10'd908: output_8x = -15757;
    10'd909: output_8x = -13314;
    10'd910: output_8x = -9305;
    10'd911: output_8x = -4382;
    10'd912: output_8x = 729;
    10'd913: output_8x = 5337;
    10'd914: output_8x = 8873;
    10'd915: output_8x = 10953;
    10'd916: output_8x = 11419;
    10'd917: output_8x = 10341;
    10'd918: output_8x = 7987;
    10'd919: output_8x = 4773;
    10'd920: output_8x = 1197;
    10'd921: output_8x = -2238;
    10'd922: output_8x = -5091;
    10'd923: output_8x = -7033;
    10'd924: output_8x = -7884;
    10'd925: output_8x = -7623;
    10'd926: output_8x = -6381;
    10'd927: output_8x = -4406;
    10'd928: output_8x = -2023;
    10'd929: output_8x = 417;
    10'd930: output_8x = 2589;
    10'd931: output_8x = 4228;
    10'd932: output_8x = 5165;
    10'd933: output_8x = 5338;
    10'd934: output_8x = 4794;
    10'd935: output_8x = 3670;
    10'd936: output_8x = 2165;
    10'd937: output_8x = 514;
    10'd938: output_8x = -1049;
    10'd939: output_8x = -2331;
    10'd940: output_8x = -3186;
    10'd941: output_8x = -3542;
    10'd942: output_8x = -3399;
    10'd943: output_8x = -2824;
    10'd944: output_8x = -1934;
    10'd945: output_8x = -877;
    10'd946: output_8x = 190;
    10'd947: output_8x = 1128;
    10'd948: output_8x = 1826;
    10'd949: output_8x = 2214;
    10'd950: output_8x = 2273;
    10'd951: output_8x = 2028;
    10'd952: output_8x = 1543;
    10'd953: output_8x = 906;
    10'd954: output_8x = 216;
    10'd955: output_8x = -427;
    10'd956: output_8x = -948;
    10'd957: output_8x = -1290;
    10'd958: output_8x = -1427;
    10'd959: output_8x = -1362;
    10'd960: output_8x = -1126;
    10'd961: output_8x = -770;
    10'd962: output_8x = -352;
    10'd963: output_8x = 63;
    10'd964: output_8x = 424;
    10'd965: output_8x = 690;
    10'd966: output_8x = 834;
    10'd967: output_8x = 853;
    10'd968: output_8x = 758;
    10'd969: output_8x = 576;
    10'd970: output_8x = 342;
    10'd971: output_8x = 90;
    10'd972: output_8x = -141;
    10'd973: output_8x = -326;
    10'd974: output_8x = -446;
    10'd975: output_8x = -493;
    10'd976: output_8x = -469;
    10'd977: output_8x = -387;
    10'd978: output_8x = -267;
    10'd979: output_8x = -126;
    10'd980: output_8x = 9;
    10'd981: output_8x = 127;
    10'd982: output_8x = 213;
    10'd983: output_8x = 259;
    10'd984: output_8x = 265;
    10'd985: output_8x = 236;
    10'd986: output_8x = 181;
    10'd987: output_8x = 110;
    10'd988: output_8x = 36;
    10'd989: output_8x = -30;
    10'd990: output_8x = -83;
    10'd991: output_8x = -117;
    10'd992: output_8x = -131;
    10'd993: output_8x = -125;
    10'd994: output_8x = -104;
    10'd995: output_8x = -72;
    10'd996: output_8x = -36;
    10'd997: output_8x = -1;
    10'd998: output_8x = 27;
    10'd999: output_8x = 47;
    10'd1000: output_8x = 59;
    10'd1001: output_8x = 62;
    10'd1002: output_8x = 55;
    10'd1003: output_8x = 45;
    10'd1004: output_8x = 30;
    10'd1005: output_8x = 16;
    10'd1006: output_8x = 2;
    10'd1007: output_8x = -7;
    10'd1008: output_8x = -13;
    10'd1009: output_8x = -17;
    10'd1010: output_8x = -16;
    10'd1011: output_8x = -14;
    10'd1012: output_8x = -19;
    default: output_8x = 0;
    endcase
    end

endmodule

